/*
* Filename:    usb_host.sv
*
* Created by:  William Cunningham
* E-mail:      wrcunnin@purdue.edu
* Date:        09/03/2025
* Description: Top level module for the USB Host
*/

module usb_host ();

endmodule
